entity Hola_Mundo is
end entity;
 
architecture sim of Hola_Mundo is
begin
 
    process is
    begin
 
        report "Hola Mundo con VHDL!";
        wait;
 
    end process;
 
end architecture;